module top_module ( input a, input b, output out );
    mod_a (a,b,out);
endmodule

